module uart_tx(

input wire sys_clk,
input wire sys_rst_n,
input wire [7:0]in_data,
input wire tx_statr_flag,

output reg tx

);

reg [31:0]rx_cnt;
reg [3:0]rx_bit_cnt;
reg bit_flag;
reg en;


localparam  CLK_FREQ = 32'd25_000_000;            // 系统时钟频率
//localparam  UART_BPS = 32'd208333;               // 串口波特率
localparam  UART_BPS = 32'd921600;               // 串口波特率
localparam  BPS_CNT  = CLK_FREQ/UART_BPS;   // 为得到指定波特率，对系统时钟计数BPS_CNT次



always @(posedge sys_clk or negedge sys_rst_n)
			if(sys_rst_n == 1'b0)
				en <= 1'b0;
			else if(tx_statr_flag == 1'b1)
				en <= 1'b1;
			else if(bit_flag == 1'b1 && rx_bit_cnt == 4'd10)
				en <= 1'b0;
			else
				en <= en;

always @(posedge sys_clk or negedge sys_rst_n)
			if(sys_rst_n == 1'b0)
				rx_cnt <= 32'd0;
			else if(rx_cnt == BPS_CNT)
				rx_cnt <= 32'd0;
			else if(en == 1'b1)
				rx_cnt <= rx_cnt + 32'd1;
			else
				rx_cnt <= 32'd0;
				
always @(posedge sys_clk or negedge sys_rst_n)
			if(sys_rst_n == 1'b0)
				bit_flag <= 1'b0;
			else if(rx_cnt == BPS_CNT >> 1)
				bit_flag <= 1'b1;
			else
				bit_flag <= 1'b0;

				
always @(posedge sys_clk or negedge sys_rst_n)
			if(sys_rst_n == 1'b0)
				rx_bit_cnt <= 4'd1;
			else if(rx_bit_cnt == 4'd10 && bit_flag == 1'b1)
				rx_bit_cnt <= 4'd1;
			else if(bit_flag == 1'b1)
				rx_bit_cnt <= rx_bit_cnt + 4'd1;
			else
				rx_bit_cnt <= rx_bit_cnt;


always @(posedge sys_clk or negedge sys_rst_n)
			if(sys_rst_n == 1'b0)
				tx <= 1'b1;
			else if(bit_flag == 1'b1)
				case (rx_bit_cnt)
					4'd1 : tx <= 1'b0;
					4'd2 : tx <= in_data[0];
					4'd3 : tx <= in_data[1];
					4'd4 : tx <= in_data[2];
					4'd5 : tx <= in_data[3];
					4'd6 : tx <= in_data[4];
					4'd7 : tx <= in_data[5];
					4'd8 : tx <= in_data[6];
					4'd9 : tx <= in_data[7];
					4'd10 : tx <= 1'b1;
					default : tx <= 1'b1;
				endcase	

endmodule
